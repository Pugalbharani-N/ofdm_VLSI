module tb_inverse_cyclic_prefix();

    // Testbench signals
    reg [303:0] symbol_out;
    wire [127:0] I_FFT;
    wire [127:0] Q_FFT;
    
    // Instantiate the module
    inverse_cyclic_prefix uut (
        .symbol_out(symbol_out),
        .I_FFT(I_FFT),
        .Q_FFT(Q_FFT)
    );

    // Test vector array (16 values)
    reg [303:0] test_vectors [0:15];
    integer i;

    initial begin
        // Initialize test vectors
        test_vectors[0]  = 304'h001400140014000a000a000a000a000a000a000a000a00140014001400140014001400140014;
        test_vectors[1]  = 304'h0014001400140005000500050005000500050005000500140014001400140014001400140014;
        test_vectors[2]  = 304'h0014001400140014001400140014001400140014001400140014001400140014001400140014;
        test_vectors[3]  = 304'h001400140014000f000f000f000f000f000f000f000f00140014001400140014001400140014;
        test_vectors[4]  = 304'h000f000f000f000a000a000a000a000a000a000a000a000f000f000f000f000f000f000f000f;
        test_vectors[5]  = 304'h000f000f000f00050005000500050005000500050005000f000f000f000f000f000f000f000f;
        test_vectors[6]  = 304'h000f000f000f00140014001400140014001400140014000f000f000f000f000f000f000f000f;
        test_vectors[7]  = 304'h000f000f000f000f000f000f000f000f000f000f000f000f000f000f000f000f000f000f000f;
        test_vectors[8]  = 304'h000a000a000a000a000a000a000a000a000a000a000a000a000a000a000a000a000a000a000a;
        test_vectors[9]  = 304'h000a000a000a00050005000500050005000500050005000a000a000a000a000a000a000a000a;
        test_vectors[10] = 304'h000a000a000a00140014001400140014001400140014000a000a000a000a000a000a000a000a;
        test_vectors[11] = 304'h000a000a000a000f000f000f000f000f000f000f000f000a000a000a000a000a000a000a000a;
        test_vectors[12] = 304'h000500050005000a000a000a000a000a000a000a000a00050005000500050005000500050005;
        test_vectors[13] = 304'h0005000500050005000500050005000500050005000500050005000500050005000500050005;
        test_vectors[14] = 304'h0005000500050014001400140014001400140014001400050005000500050005000500050005;
        test_vectors[15] = 304'h000500050005000f000f000f000f000f000f000f000f00050005000500050005000500050005;

        // Apply each test vector
        for (i = 0; i < 16; i = i + 1) begin
            symbol_out = test_vectors[i];
            #10; // Wait for processing
            $display("Test %0d: I_FFT = %h, Q_FFT = %h", i, I_FFT, Q_FFT);
        end

        // Finish simulation
        $finish;
    end

endmodule


